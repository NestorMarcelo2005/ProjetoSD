// Verilog test fixture created from schematic C:\Users\nESTOR\Desktop\trabalhos\Balanca\projetof.sch - Fri Nov 10 14:18:14 2023

`timescale 1ns / 1ps

module projetof_projetof_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   projetof UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
